module hilo_reg
(
    
)

endmodule