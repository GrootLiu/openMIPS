/*
 * @Author: Groot
 * @Date: 2022-04-13 16:14:33
 * @LastEditTime: 2022-04-14 15:14:19
 * @LastEditors: Groot
 * @Description: 
 * @FilePath: /openMIPS/vsrc/hilo_reg.v
 * 版权声明
 */
`include "./include/define.v"

module hilo_reg
(
    
)

endmodule