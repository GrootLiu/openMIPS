/*
 * @Author: Groot
 * @Date: 2022-04-09 18:01:23
 * @LastEditTime: 2022-04-14 15:41:39
 * @LastEditors: Groot
 * @Description:
 * @FilePath: /openMIPS/vsrc/id_ex.v
 * 版权声明
 */
`include "/home/groot/openMIPS/include/define.v"

module id_ex (input wire clk,
              input wire rst,
              input wire[`AluOpBus] id_aluop,
              input wire [`AluSelBus] id_alusel,
              input wire[`RegBus] id_reg1,
              input wire[`RegBus] id_reg2,
              input wire[`RegAddBus] id_wd,
              input wire id_wreg,
              output reg[`AluOpBus] ex_aluop,
              output reg[`AluSelBus] ex_alusel,
              output reg[`RegBus] ex_reg1,
              output reg[`RegBus] ex_reg2,
              output reg[`RegAddBus] ex_wd,
              output reg ex_wreg);
    
    always @(posedge clk)
    begin
        if (rst == `RstEnable)
        begin
            ex_aluop  <= `EXE_NOP_OP;
            ex_alusel <= `EXE_RES_NOP;
            ex_reg1   <= `ZeroWord;
            ex_reg2   <= `ZeroWord;
            ex_wd     <= `NOPRegAddr;
            ex_wreg   <= `WriteDisable;
        end
        else
        begin
            ex_aluop  <= id_aluop;
            ex_alusel <= id_alusel;
            ex_reg1   <= id_reg1;
            ex_reg2   <= id_reg2;
            ex_wd     <= id_wd;
            ex_wreg   <= id_wreg;
        end
    end
    
endmodule //id_ex
